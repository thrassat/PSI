`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:17:37 05/10/2019 
// Design Name: 
// Module Name:    banc_registre 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module banc_registre(
    input [3:0] aA,
    input [3:0] aB,
    input [3:0] aW,
    input W,
    input [7:0] DATA,
    input RST,
    input CLK,
    output [7:0] QA,
    output [7:0] QB
    );


endmodule
