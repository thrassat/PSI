----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:21:45 05/13/2019 
-- Design Name: 
-- Module Name:    mux - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mux is
	 generic (N:natural := 16) ; 
    Port ( i0 : in  STD_LOGIC_VECTOR (N-1 downto 0);
           i1 : in  STD_LOGIC_VECTOR (N-1 downto 0);
           sel : in  STD_LOGIC ; 
           S : out  STD_LOGIC_VECTOR (N-1 downto 0));
end mux;

architecture Behavioral of mux is

begin
	S <= i0 WHEN sel='0' else 
		  i1 ; 


end Behavioral;

